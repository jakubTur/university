CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 120 30 120 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 298 272 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -19 8 -11
1 D
-3 -32 4 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 421 309 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-6 -25 1 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 429 254 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -17 7 -9
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 423 203 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
5 4011~
219 348 271 0 3 22
0 10 10 3
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 5 0
1 U
5394 0 0
0
0
5 4011~
219 491 305 0 3 22
0 12 12 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 5 0
1 U
7734 0 0
0
0
5 4011~
219 491 254 0 3 22
0 13 13 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 5 0
1 U
9914 0 0
0
0
5 4011~
219 490 203 0 3 22
0 14 14 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3747 0 0
0
0
9 2-In AND~
219 429 414 0 3 22
0 11 3 4
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1743344971
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
7 Ground~
168 622 418 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 584 407 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
14 Logic Display~
6 562 458 0 1 2
10 15
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
7 74LS151
20 484 435 0 14 29
0 16 17 18 19 4 4 4 3 2
2 13 14 15 20
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
14 Logic Display~
6 741 257 0 1 2
10 6
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
5 4023~
219 596 225 0 4 22
0 9 3 8 5
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
7668 0 0
0
0
5 4011~
219 686 261 0 3 22
0 5 7 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
4718 0 0
0
0
5 4011~
219 605 314 0 3 22
0 11 3 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3874 0 0
0
0
27
0 8 3 0 0 8192 0 0 13 14 0 4
375 323
376 323
376 471
452 471
0 7 4 0 0 8320 0 0 13 3 0 3
427 444
427 462
452 462
0 6 4 0 0 0 0 0 13 4 0 4
427 444
444 444
444 453
452 453
3 5 4 0 0 0 0 9 13 0 0 3
427 437
427 444
452 444
4 1 5 0 0 4224 0 15 16 0 0 4
623 225
654 225
654 252
662 252
3 1 6 0 0 4224 0 16 14 0 0 2
713 261
725 261
3 2 7 0 0 8320 0 17 16 0 0 4
632 314
654 314
654 270
662 270
3 2 3 0 0 12288 0 5 15 0 0 4
375 271
376 271
376 225
572 225
3 3 8 0 0 4224 0 7 15 0 0 4
518 254
564 254
564 234
572 234
3 1 9 0 0 4224 0 8 15 0 0 4
517 203
564 203
564 216
572 216
2 0 3 0 0 0 0 9 0 0 14 2
418 392
418 323
2 1 10 0 0 12288 0 5 1 0 0 4
324 280
319 280
319 272
310 272
1 1 10 0 0 8320 0 5 1 0 0 4
324 262
319 262
319 272
310 272
3 2 3 0 0 8320 0 5 17 0 0 3
375 271
375 323
581 323
0 1 11 0 0 8320 0 0 9 16 0 4
532 305
532 338
436 338
436 392
3 1 11 0 0 0 0 6 17 0 0 2
518 305
581 305
1 2 12 0 0 4224 0 2 6 0 0 4
433 309
459 309
459 314
467 314
1 1 12 0 0 0 0 2 6 0 0 4
433 309
459 309
459 296
467 296
0 11 13 0 0 4224 0 0 13 20 0 5
454 254
454 380
530 380
530 426
516 426
1 2 13 0 0 0 0 3 7 0 0 4
441 254
459 254
459 263
467 263
1 1 13 0 0 0 0 3 7 0 0 4
441 254
459 254
459 245
467 245
0 12 14 0 0 4224 0 0 13 23 0 5
447 203
447 486
530 486
530 435
516 435
1 2 14 0 0 0 0 4 8 0 0 4
435 203
458 203
458 212
466 212
1 1 14 0 0 0 0 4 8 0 0 4
435 203
458 203
458 194
466 194
13 1 15 0 0 4224 0 13 12 0 0 2
516 462
546 462
10 1 2 0 0 4224 0 13 10 0 0 6
516 417
573 417
573 422
607 422
607 419
615 419
9 1 2 0 0 0 0 13 11 0 0 2
522 408
577 408
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1836704 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 2
1
425 205
0 0 0 0 0	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
