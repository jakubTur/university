CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 1 120 9
38 94 1498 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 94 1498 791
177209362 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 108 300 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 110 238 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 109 154 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
5 SCOPE
12 89 72 0 1 11
0 3
0
0 0 57584 0
1 B
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 126 74 0 1 11
0 4
0
0 0 57584 0
1 C
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 54 72 0 1 11
0 5
0
0 0 57584 0
1 A
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 495 186 0 1 11
0 6
0
0 0 57584 0
1 F
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 4011~
219 364 230 0 3 22
0 3 9 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3747 0 0
0
0
5 4011~
219 364 188 0 3 22
0 8 5 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3549 0 0
0
0
5 4011~
219 156 262 0 3 22
0 4 4 13
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
7931 0 0
0
0
5 4011~
219 154 189 0 3 22
0 3 3 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
9325 0 0
0
0
5 4011~
219 171 133 0 3 22
0 5 5 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
8903 0 0
0
0
7 Ground~
168 350 401 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 306 385 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
8 2-In OR~
219 25 384 0 3 22
0 3 5 14
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
7668 0 0
0
0
8 2-In OR~
219 80 382 0 3 22
0 9 8 15
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1809612885
65 0 0 0 4 1 5 0
1 U
4718 0 0
0
0
14 Logic Display~
6 274 427 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
7 Ground~
168 266 376 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 74LS151
20 173 404 0 14 29
0 17 18 19 20 21 22 14 15 2
2 2 4 16 23
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
14 Logic Display~
6 534 210 0 1 2
10 6
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
5 4012~
219 451 214 0 5 22
0 7 11 10 12 6
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 -1810453831
65 0 0 0 2 1 4 0
1 U
3750 0 0
0
0
5 4011~
219 363 291 0 3 22
0 5 4 12
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
8778 0 0
0
0
5 4011~
219 360 142 0 3 22
0 9 13 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1642681677
65 0 0 0 4 1 1 0
1 U
538 0 0
0
0
34
1 0 3 0 0 4096 0 4 0 0 19 2
89 84
89 198
1 0 4 0 0 4096 0 5 0 0 33 4
126 86
126 295
136 295
136 300
1 0 5 0 0 4096 0 6 0 0 22 2
54 84
54 129
1 0 6 0 0 4096 0 7 0 0 32 2
495 198
495 214
3 1 7 0 0 8320 0 23 21 0 0 4
387 142
419 142
419 201
427 201
0 2 8 0 0 4096 0 0 16 9 0 4
201 189
201 330
74 330
74 366
0 1 3 0 0 4224 0 0 8 19 0 2
122 221
340 221
2 0 9 0 0 8192 0 8 0 0 21 3
340 239
241 239
241 133
3 1 8 0 0 4224 0 11 9 0 0 4
181 189
332 189
332 179
340 179
0 2 5 0 0 0 0 0 9 34 0 3
302 166
302 197
340 197
3 3 10 0 0 8320 0 8 21 0 0 3
391 230
391 219
427 219
3 2 11 0 0 8320 0 9 21 0 0 3
391 188
391 210
427 210
3 4 12 0 0 8320 0 22 21 0 0 4
390 291
419 291
419 228
427 228
3 2 13 0 0 8320 0 10 23 0 0 3
183 262
183 151
336 151
1 2 4 0 0 0 0 1 10 0 0 4
120 300
126 300
126 271
132 271
1 1 4 0 0 0 0 1 10 0 0 4
120 300
126 300
126 253
132 253
0 2 3 0 0 0 0 0 11 19 0 3
122 202
122 198
130 198
0 1 3 0 0 0 0 0 11 19 0 3
122 198
122 180
130 180
1 1 3 0 0 0 0 2 15 0 0 4
122 238
122 198
37 198
37 368
0 1 9 0 0 4224 0 0 16 21 0 4
213 133
213 349
92 349
92 366
3 1 9 0 0 0 0 12 23 0 0 2
198 133
336 133
1 2 5 0 0 12416 0 3 15 0 0 4
121 154
121 129
19 129
19 368
1 1 5 0 0 0 0 3 12 0 0 4
121 154
141 154
141 124
147 124
1 2 5 0 0 0 0 3 12 0 0 4
121 154
141 154
141 142
147 142
11 1 2 0 0 4224 0 19 13 0 0 4
205 395
295 395
295 402
343 402
10 1 2 0 0 0 0 19 14 0 0 6
205 386
255 386
255 391
291 391
291 386
299 386
3 7 14 0 0 8320 0 15 19 0 0 3
28 414
28 431
141 431
3 8 15 0 0 8320 0 16 19 0 0 3
83 412
83 440
141 440
13 1 16 0 0 4224 0 19 17 0 0 2
205 431
258 431
9 1 2 0 0 0 0 19 18 0 0 2
211 377
259 377
12 0 4 0 0 0 0 19 0 0 33 3
205 404
236 404
236 300
5 1 6 0 0 4224 0 21 20 0 0 2
478 214
518 214
1 2 4 0 0 4224 0 1 22 0 0 2
120 300
339 300
1 1 5 0 0 0 0 3 22 0 0 5
121 154
121 166
331 166
331 282
339 282
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
