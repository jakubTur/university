CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
580 130 1 200 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 597 264 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 597 227 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-9 -16 5 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
7 Ground~
168 640 323 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 682 284 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
4 LED~
171 1292 213 0 1 2
10 4
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5394 0 0
0
0
4 LED~
171 1219 211 0 1 2
10 5
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7734 0 0
0
0
4 LED~
171 1103 206 0 1 2
10 6
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9914 0 0
0
0
4 LED~
171 1030 204 0 1 2
10 7
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3747 0 0
0
0
10 3-In NAND~
219 879 315 0 4 22
0 4 5 6 8
0
0 0 624 270
6 74LS10
-21 -28 21 -20
3 U2A
19 -7 40 1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
3549 0 0
0
0
7 74LS194
49 772 262 0 14 29
0 9 3 2 2 8 3 10 11 12
13 4 5 6 7
0
0 0 13040 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
13
4 1 2 0 0 4224 0 10 3 0 0 3
740 271
640 271
640 317
1 0 3 0 0 4224 0 1 0 0 12 4
609 264
721 264
721 265
726 265
0 1 4 0 0 8320 0 0 5 10 0 4
889 271
889 200
1292 200
1292 203
0 1 5 0 0 8320 0 0 6 9 0 4
880 280
880 195
1219 195
1219 201
0 1 6 0 0 8320 0 0 7 8 0 5
871 282
871 190
1100 190
1100 196
1103 196
14 1 7 0 0 12416 0 10 8 0 0 5
804 298
861 298
861 186
1030 186
1030 194
1 3 2 0 0 0 0 4 10 0 0 3
682 278
682 253
740 253
13 3 6 0 0 0 0 10 9 0 0 5
804 289
861 289
861 282
871 282
871 290
12 2 5 0 0 0 0 10 9 0 0 3
804 280
880 280
880 290
11 1 4 0 0 0 0 10 9 0 0 3
804 271
889 271
889 290
5 4 8 0 0 12416 0 10 9 0 0 5
740 280
730 280
730 349
880 349
880 341
2 6 3 0 0 0 0 10 10 0 0 4
740 244
726 244
726 298
734 298
1 1 9 0 0 8320 0 2 10 0 0 3
609 227
609 226
740 226
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1246186 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 100 100 0 0
77 66 1487 276
0 0 0 0
1487 66
77 66
1487 66
1487 276
0 0
9.99575e-007 0 4.57143 4.14286 1e-006 1e-006
12409 0
0 3e-007 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
