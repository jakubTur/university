CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 120 1 100 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 816
177209362 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 691 482 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 501 598 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 769 297 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 975 166 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 410 172 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 204 303 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
9 Inverter~
13 687 626 0 2 22
0 3 5
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4E
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 4 0
1 U
9914 0 0
0
0
9 Inverter~
13 556 599 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 4 0
1 U
3747 0 0
0
0
9 2-In AND~
219 675 599 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 9 0
1 U
3549 0 0
0
0
14 Logic Display~
6 1000 616 0 1 2
10 10
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 Z1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 870 628 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 863 517 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
9 2-In AND~
219 948 620 0 3 22
0 8 11 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 9 0
1 U
3834 0 0
0
0
7 Ground~
168 740 749 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
5 4027~
219 790 697 0 7 32
0 2 8 3 6 4 9 11
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 2 5 0
1 U
7668 0 0
0
0
5 4027~
219 790 587 0 7 32
0 2 7 3 9 4 38 8
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5A
20 -57 41 -49
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 1390027930
65 0 0 512 2 1 5 0
1 U
4718 0 0
0
0
10 2-In NAND~
219 1152 288 0 3 22
0 13 12 15
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 8 0
1 U
3874 0 0
0
0
10 2-In NAND~
219 927 370 0 3 22
0 19 18 17
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 8 0
1 U
6671 0 0
0
0
10 2-In NAND~
219 930 286 0 3 22
0 20 19 16
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 7 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 842 379 0 3 22
0 21 13 18
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 7 0
1 U
4871 0 0
0
0
10 2-In NAND~
219 842 326 0 3 22
0 21 12 19
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 7 0
1 U
3750 0 0
0
0
10 2-In NAND~
219 842 252 0 3 22
0 22 21 20
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 1574577301
65 0 0 0 4 1 7 0
1 U
8778 0 0
0
0
5 4013~
219 1051 313 0 6 22
0 2 16 23 2 22 13
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 2 6 0
1 U
538 0 0
0
0
5 4013~
219 1054 401 0 6 22
0 2 17 23 2 39 12
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 6 0
1 U
6843 0 0
0
0
9 Inverter~
13 1205 287 0 2 22
0 15 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 4 0
1 U
3136 0 0
0
0
7 Ground~
168 1022 466 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
14 Logic Display~
6 1255 282 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
1 Z
-2 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 1100 228 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 1200 343 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 635 349 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
14 Logic Display~
6 537 236 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
14 Logic Display~
6 638 288 0 1 2
10 27
0
0 0 53872 270
6 100MEG
3 -16 45 -8
1 Z
-2 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4551 0 0
0
0
7 Ground~
168 457 472 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3635 0 0
0
0
9 Inverter~
13 551 349 0 2 22
0 28 29
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
3973 0 0
0
0
9 Inverter~
13 373 332 0 2 22
0 28 32
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
3851 0 0
0
0
8 2-In OR~
219 368 373 0 3 22
0 36 35 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
8383 0 0
0
0
8 2-In OR~
219 371 283 0 3 22
0 30 36 34
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2062367692
65 0 0 0 4 1 3 0
1 U
9334 0 0
0
0
9 2-In AND~
219 585 292 0 3 22
0 25 29 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
7471 0 0
0
0
9 2-In AND~
219 279 382 0 3 22
0 37 25 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3334 0 0
0
0
9 2-In AND~
219 280 312 0 3 22
0 37 32 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3559 0 0
0
0
9 2-In AND~
219 280 274 0 3 22
0 31 37 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1961704390
65 0 0 0 4 1 2 0
1 U
984 0 0
0
0
5 4013~
219 489 407 0 6 22
0 2 33 24 2 28 26
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 2 1 0
1 U
7557 0 0
0
0
5 4013~
219 486 319 0 6 22
0 2 34 24 2 31 25
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 1 0
1 U
3146 0 0
0
0
68
1 0 3 0 0 8192 0 7 0 0 18 3
708 626
708 625
726 625
3 5 4 0 0 8320 0 9 15 0 0 5
696 599
761 599
761 711
790 711
790 703
3 5 4 0 0 0 0 9 16 0 0 3
696 599
790 599
790 593
0 1 2 0 0 4096 0 0 15 5 0 3
740 632
790 632
790 640
1 1 2 0 0 12416 0 16 14 0 0 4
790 530
790 526
740 526
740 743
2 2 5 0 0 8320 0 9 7 0 0 4
651 608
651 625
672 625
672 626
0 1 6 0 0 8192 0 0 9 9 0 3
626 599
626 590
651 590
1 2 7 0 0 12416 0 2 16 0 0 4
513 598
537 598
537 551
766 551
2 4 6 0 0 12416 0 8 15 0 0 4
577 599
626 599
626 679
766 679
1 1 7 0 0 0 0 2 8 0 0 4
513 598
533 598
533 599
541 599
0 2 8 0 0 8192 0 0 15 17 0 5
841 551
841 615
758 615
758 661
766 661
6 4 9 0 0 8320 0 15 16 0 0 6
820 679
824 679
824 512
758 512
758 569
766 569
3 1 10 0 0 4224 0 13 10 0 0 2
969 620
984 620
1 0 11 0 0 4096 0 11 0 0 16 2
870 646
870 661
1 0 8 0 0 0 0 12 0 0 17 2
863 535
863 551
7 2 11 0 0 4224 0 15 13 0 0 4
814 661
916 661
916 629
924 629
7 1 8 0 0 4224 0 16 13 0 0 4
814 551
916 551
916 611
924 611
0 3 3 0 0 4224 0 0 15 19 0 3
726 560
726 670
766 670
3 1 3 0 0 0 0 16 1 0 0 4
766 560
726 560
726 482
703 482
2 0 12 0 0 8192 0 17 0 0 39 3
1128 297
1124 297
1124 365
0 1 13 0 0 4096 0 0 17 31 0 5
1079 277
1079 323
1120 323
1120 279
1128 279
2 1 14 0 0 12416 0 25 27 0 0 4
1226 287
1232 287
1232 286
1239 286
3 1 15 0 0 12416 0 17 25 0 0 4
1179 288
1184 288
1184 287
1190 287
3 2 16 0 0 4224 0 19 23 0 0 4
957 286
1019 286
1019 277
1027 277
3 2 17 0 0 4224 0 18 24 0 0 4
954 370
1022 370
1022 365
1030 365
2 3 18 0 0 4224 0 18 20 0 0 2
903 379
869 379
3 1 19 0 0 8320 0 21 18 0 0 4
869 326
895 326
895 361
903 361
2 3 19 0 0 0 0 19 21 0 0 4
906 295
895 295
895 326
869 326
3 1 20 0 0 4224 0 22 19 0 0 4
869 252
898 252
898 277
906 277
1 1 21 0 0 8320 0 3 20 0 0 4
781 297
802 297
802 370
818 370
6 2 13 0 0 12416 0 23 20 0 0 6
1075 277
1095 277
1095 412
810 412
810 388
818 388
6 2 12 0 0 12416 0 24 21 0 0 8
1078 365
1088 365
1088 335
873 335
873 346
810 346
810 335
818 335
1 1 21 0 0 0 0 3 21 0 0 4
781 297
803 297
803 317
818 317
1 2 21 0 0 0 0 3 22 0 0 4
781 297
802 297
802 261
818 261
5 1 22 0 0 12416 0 23 22 0 0 6
1081 295
1085 295
1085 232
810 232
810 243
818 243
0 3 23 0 0 8192 0 0 24 37 0 5
984 295
985 295
985 384
1030 384
1030 383
1 3 23 0 0 8320 0 4 23 0 0 4
987 166
984 166
984 295
1027 295
0 1 13 0 0 0 0 0 28 21 0 2
1100 323
1100 246
6 1 12 0 0 0 0 24 29 0 0 3
1078 365
1200 365
1200 361
4 0 2 0 0 0 0 24 0 0 43 3
1054 407
1054 405
1022 405
1 0 2 0 0 0 0 24 0 0 43 3
1054 344
1054 340
1022 340
4 0 2 0 0 0 0 23 0 0 43 3
1051 319
1051 323
1022 323
1 1 2 0 0 128 0 23 26 0 0 4
1051 256
1051 252
1022 252
1022 460
0 3 24 0 0 8192 0 0 42 45 0 4
454 301
457 301
457 389
465 389
1 3 24 0 0 8320 0 5 43 0 0 4
422 172
454 172
454 301
462 301
0 1 25 0 0 4096 0 0 31 58 0 2
537 283
537 254
6 1 26 0 0 4224 0 42 30 0 0 3
513 371
635 371
635 367
3 1 27 0 0 4224 0 38 32 0 0 2
606 292
622 292
4 0 2 0 0 0 0 42 0 0 52 3
489 413
489 411
457 411
1 0 2 0 0 0 0 42 0 0 52 3
489 350
489 346
457 346
4 0 2 0 0 0 0 43 0 0 52 3
486 325
486 329
457 329
1 1 2 0 0 0 0 43 33 0 0 4
486 262
486 258
457 258
457 466
0 2 25 0 0 8320 0 0 39 58 0 5
539 283
539 418
247 418
247 391
255 391
1 5 28 0 0 12288 0 34 42 0 0 4
554 367
553 367
553 389
519 389
2 2 29 0 0 8320 0 38 34 0 0 4
561 301
553 301
553 331
554 331
3 1 30 0 0 4224 0 41 37 0 0 2
301 274
358 274
5 1 31 0 0 12416 0 43 41 0 0 6
516 301
520 301
520 240
247 240
247 265
256 265
6 1 25 0 0 0 0 43 38 0 0 2
510 283
561 283
1 5 28 0 0 4224 0 35 42 0 0 4
394 332
523 332
523 389
519 389
2 2 32 0 0 12416 0 40 35 0 0 4
256 321
248 321
248 332
358 332
3 2 33 0 0 4224 0 36 42 0 0 4
401 373
457 373
457 371
465 371
3 2 34 0 0 4224 0 37 43 0 0 2
404 283
462 283
3 2 35 0 0 4224 0 39 36 0 0 2
300 382
355 382
3 1 36 0 0 8192 0 40 36 0 0 3
301 312
301 364
355 364
3 2 36 0 0 8320 0 40 37 0 0 3
301 312
301 292
358 292
1 1 37 0 0 4096 0 6 40 0 0 2
216 303
256 303
1 1 37 0 0 4224 0 6 39 0 0 3
216 303
216 373
255 373
1 2 37 0 0 0 0 6 41 0 0 3
216 303
216 283
256 283
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1181174 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 2 2
1
205 303
0 0 0 0 0	6 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
