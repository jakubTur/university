CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 260 1 120 9
38 95 1498 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 703 1498 791
193986578 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 92 369 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 145 370 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 203 372 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 251 372 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
5 SCOPE
12 731 520 0 1 11
0 3
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 565 532 0 1 11
0 4
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
14 Logic Display~
6 533 579 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
5 4013~
219 659 576 0 6 22
0 2 5 4 2 5 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 3 0
1 U
3747 0 0
0
0
14 Logic Display~
6 765 536 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
7 Ground~
168 659 600 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 636 482 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
5 4023~
219 354 501 0 4 22
0 10 6 11 12
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 8 0
1 U
8903 0 0
0
0
9 Inverter~
13 171 420 0 2 22
0 8 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 512 6 6 5 0
1 U
3834 0 0
0
0
9 Inverter~
13 109 420 0 2 22
0 15 10
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 5 0
1 U
3363 0 0
0
0
9 Inverter~
13 226 421 0 2 22
0 9 11
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 5 0
1 U
7668 0 0
0
0
9 Inverter~
13 276 420 0 2 22
0 7 6
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 5 0
1 U
4718 0 0
0
0
5 4023~
219 354 554 0 4 22
0 10 8 7 14
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 8 0
1 U
3874 0 0
0
0
5 4023~
219 353 611 0 4 22
0 9 8 7 13
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 6 0
1 U
6671 0 0
0
0
5 4023~
219 450 554 0 4 22
0 12 14 13 4
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 6 0
1 U
3789 0 0
0
0
24
1 0 3 0 0 4096 0 5 0 0 7 3
731 532
731 540
730 540
1 0 4 0 0 4096 0 6 0 0 4 3
565 544
565 554
563 554
1 0 4 0 0 8192 0 7 0 0 4 3
517 583
514 583
514 554
4 3 4 0 0 4224 0 19 8 0 0 4
477 554
627 554
627 558
635 558
1 4 2 0 0 4096 0 10 8 0 0 2
659 594
659 582
1 1 2 0 0 12416 0 11 8 0 0 4
636 476
636 472
659 472
659 519
6 1 3 0 0 4224 0 8 9 0 0 2
683 540
749 540
5 2 5 0 0 12416 0 8 8 0 0 6
689 558
693 558
693 514
627 514
627 540
635 540
2 2 6 0 0 4224 0 16 12 0 0 3
279 438
279 501
330 501
0 3 7 0 0 8192 0 0 18 13 0 3
251 563
251 620
329 620
0 2 8 0 0 8192 0 0 18 14 0 3
145 554
145 611
329 611
0 1 9 0 0 4224 0 0 18 22 0 3
203 395
203 602
329 602
0 3 7 0 0 4224 0 0 17 21 0 3
251 390
251 563
330 563
0 2 8 0 0 8320 0 0 17 23 0 3
145 394
145 554
330 554
0 1 10 0 0 8320 0 0 17 17 0 3
112 492
112 545
330 545
2 3 11 0 0 8320 0 15 12 0 0 3
229 439
229 510
330 510
2 1 10 0 0 0 0 14 12 0 0 3
112 438
112 492
330 492
1 4 12 0 0 8320 0 19 12 0 0 4
426 545
389 545
389 501
381 501
4 3 13 0 0 8320 0 18 19 0 0 4
380 611
424 611
424 563
426 563
4 2 14 0 0 4224 0 17 19 0 0 2
381 554
426 554
1 1 7 0 0 0 0 4 16 0 0 4
251 384
251 397
279 397
279 402
1 1 9 0 0 0 0 3 15 0 0 4
203 384
203 395
229 395
229 403
1 1 8 0 0 0 0 2 13 0 0 4
145 382
145 394
174 394
174 402
1 1 15 0 0 8320 0 1 14 0 0 4
92 381
92 394
112 394
112 402
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
