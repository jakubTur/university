CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 30 1 200 9
38 95 1498 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 703 1498 791
193986578 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 227 79 0 1 11
0 21
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 179 79 0 1 11
0 22
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 121 77 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 68 76 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
5 SCOPE
12 623 228 0 1 11
0 3
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 493 247 0 1 11
0 4
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
7 Ground~
168 547 195 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 570 313 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
14 Logic Display~
6 650 243 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
5 4013~
219 570 283 0 6 22
0 2 5 4 2 5 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 6 0
1 U
7931 0 0
0
0
14 Logic Display~
6 473 319 0 1 2
10 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
5 4012~
219 422 265 0 5 22
0 17 16 15 14 4
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 -568416708
65 0 0 0 2 1 4 0
1 U
8903 0 0
0
0
5 4023~
219 328 376 0 4 22
0 18 19 20 14
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 3 0
1 U
3834 0 0
0
0
5 4023~
219 329 318 0 4 22
0 22 18 21 15
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 1 0
1 U
3363 0 0
0
0
5 4023~
219 330 261 0 4 22
0 20 18 21 16
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 1 0
1 U
7668 0 0
0
0
9 Inverter~
13 252 127 0 2 22
0 21 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 2 0
1 U
4718 0 0
0
0
9 Inverter~
13 202 128 0 2 22
0 22 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 2 0
1 U
3874 0 0
0
0
9 Inverter~
13 85 127 0 2 22
0 23 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
6671 0 0
0
0
9 Inverter~
13 147 127 0 2 22
0 18 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 512 6 1 2 0
1 U
3789 0 0
0
0
5 4023~
219 330 208 0 4 22
0 20 13 19 17
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 1 0
1 U
4871 0 0
0
0
28
1 0 3 0 0 4096 0 5 0 0 5 3
623 240
623 247
624 247
1 0 4 0 0 4096 0 6 0 0 7 3
493 259
493 265
491 265
1 4 2 0 0 4096 0 8 10 0 0 2
570 307
570 289
1 1 2 0 0 12416 0 7 10 0 0 4
547 189
547 185
570 185
570 226
6 1 3 0 0 4224 0 10 9 0 0 2
594 247
634 247
5 2 5 0 0 12416 0 10 10 0 0 6
600 265
604 265
604 214
538 214
538 247
546 247
5 3 4 0 0 4224 0 12 10 0 0 2
449 265
546 265
5 1 4 0 0 0 0 12 11 0 0 3
449 265
457 265
457 323
2 2 13 0 0 4224 0 16 20 0 0 3
255 145
255 208
306 208
4 4 14 0 0 8320 0 13 12 0 0 3
355 376
398 376
398 279
4 3 15 0 0 8320 0 14 12 0 0 4
356 318
390 318
390 270
398 270
4 2 16 0 0 4224 0 15 12 0 0 2
357 261
398 261
4 1 17 0 0 8320 0 20 12 0 0 4
357 208
390 208
390 252
398 252
0 1 18 0 0 8192 0 0 13 18 0 3
124 318
124 367
304 367
0 2 19 0 0 4224 0 0 13 23 0 3
205 217
205 376
304 376
0 3 20 0 0 8192 0 0 13 22 0 3
88 251
88 385
304 385
0 3 21 0 0 8192 0 0 14 20 0 3
227 270
227 327
305 327
0 2 18 0 0 8192 0 0 14 21 0 3
121 261
121 318
305 318
0 1 22 0 0 4224 0 0 14 26 0 3
179 102
179 309
305 309
0 3 21 0 0 4224 0 0 15 25 0 3
227 97
227 270
306 270
0 2 18 0 0 8320 0 0 15 27 0 3
121 101
121 261
306 261
0 1 20 0 0 8320 0 0 15 24 0 3
88 199
88 252
306 252
2 3 19 0 0 0 0 17 20 0 0 3
205 146
205 217
306 217
2 1 20 0 0 0 0 18 20 0 0 3
88 145
88 199
306 199
1 1 21 0 0 0 0 1 16 0 0 4
227 91
227 104
255 104
255 109
1 1 22 0 0 0 0 2 17 0 0 4
179 91
179 102
205 102
205 110
1 1 18 0 0 0 0 3 19 0 0 4
121 89
121 101
150 101
150 109
1 1 23 0 0 8320 0 4 18 0 0 4
68 88
68 101
88 101
88 109
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
