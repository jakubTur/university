CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
38 95 1498 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 95 1498 791
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 120 224 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 30 127 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 444 304 0 1 2
10 8
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 Z1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 443 371 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 Z2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
9 2-In AND~
219 373 310 0 3 22
0 6 4 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
5394 0 0
0
0
9 2-In AND~
219 376 375 0 3 22
0 5 6 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 4 0
1 U
7734 0 0
0
0
7 Ground~
168 209 435 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
5 4027~
219 234 347 0 7 32
0 2 6 3 6 2 5 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 466936580
65 0 0 0 2 1 5 0
1 U
3747 0 0
0
0
9 2-In AND~
219 352 197 0 3 22
0 13 12 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3549 0 0
0
0
9 2-In AND~
219 349 132 0 3 22
0 11 14 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7931 0 0
0
0
14 Logic Display~
6 419 193 0 1 2
10 9
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 Z2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 420 126 0 1 2
10 10
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 Z1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
8 2-In OR~
219 201 107 0 3 22
0 17 16 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 450224900
65 0 0 0 4 1 3 0
1 U
3834 0 0
0
0
9 2-In AND~
219 144 91 0 3 22
0 15 11 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3363 0 0
0
0
9 2-In AND~
219 153 133 0 3 22
0 6 12 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 450224900
65 0 0 0 4 1 2 0
1 U
7668 0 0
0
0
9 Inverter~
13 79 82 0 2 22
0 6 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
4718 0 0
0
0
12 D Flip-Flop~
219 270 242 0 4 9
0 18 3 12 11
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 D2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
12 D Flip-Flop~
219 272 169 0 4 9
0 11 3 14 13
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 D1
-6 -65 8 -57
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
28
0 3 3 0 0 4096 0 0 8 27 0 3
150 224
150 320
210 320
7 2 4 0 0 4224 0 8 5 0 0 4
258 311
341 311
341 319
349 319
6 1 5 0 0 4224 0 8 6 0 0 4
264 329
344 329
344 366
352 366
0 2 6 0 0 4096 0 0 8 6 0 3
197 257
197 311
210 311
0 2 6 0 0 4096 0 0 6 6 0 3
326 257
326 384
352 384
0 1 6 0 0 8192 0 0 5 11 0 5
171 329
171 257
341 257
341 301
349 301
3 1 7 0 0 4224 0 6 4 0 0 2
397 375
427 375
3 1 8 0 0 4224 0 5 3 0 0 4
394 310
421 310
421 308
428 308
1 0 2 0 0 12416 0 8 0 0 10 4
234 290
234 266
208 266
208 397
5 1 2 0 0 0 0 8 7 0 0 6
234 353
234 397
208 397
208 397
209 397
209 429
0 4 6 0 0 4224 0 0 8 20 0 3
65 125
65 329
210 329
3 1 9 0 0 4224 0 9 11 0 0 2
373 197
403 197
3 1 10 0 0 4224 0 10 12 0 0 4
370 132
397 132
397 130
404 130
0 1 11 0 0 4096 0 0 10 28 0 2
306 123
325 123
0 2 12 0 0 8192 0 0 9 19 0 4
306 227
320 227
320 206
328 206
4 1 13 0 0 8320 0 18 9 0 0 4
296 133
320 133
320 188
328 188
3 2 14 0 0 4224 0 18 10 0 0 4
302 151
317 151
317 141
325 141
0 2 11 0 0 4224 0 0 14 28 0 4
306 181
112 181
112 100
120 100
3 2 12 0 0 12416 0 17 15 0 0 8
300 224
306 224
306 247
194 247
194 165
96 165
96 142
129 142
0 1 6 0 0 0 0 0 15 25 0 4
54 127
54 125
129 125
129 124
2 1 15 0 0 4224 0 16 14 0 0 2
100 82
120 82
2 3 16 0 0 8320 0 13 15 0 0 4
188 116
182 116
182 133
174 133
3 1 17 0 0 4224 0 14 13 0 0 4
165 91
180 91
180 98
188 98
3 1 18 0 0 8320 0 13 17 0 0 4
234 107
238 107
238 206
246 206
1 1 6 0 0 0 0 2 16 0 0 4
42 127
54 127
54 82
64 82
0 2 3 0 0 0 0 0 18 27 0 3
228 224
228 151
248 151
1 2 3 0 0 4224 0 1 17 0 0 2
132 224
246 224
4 1 11 0 0 0 0 17 18 0 0 6
294 206
306 206
306 119
240 119
240 133
248 133
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
917950 1079360 100 100 0 0
0 0 0 0
5 88 166 158
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
