CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
330 140 1 200 9
38 95 1498 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 95 1498 791
143654930 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 391 236 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 410 309 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-4 -24 10 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 519 215 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
7 Ground~
168 440 376 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 694 297 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
14 Logic Display~
6 997 261 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 929 240 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 853 212 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 767 208 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
7 74LS194
49 587 352 0 14 29
0 7 9 8 2 6 9 9 2 2
2 3 4 5 6
0
0 0 13040 0
7 74LS194
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
14
11 1 3 0 0 4224 0 10 9 0 0 3
619 361
767 361
767 226
12 1 4 0 0 4224 0 10 8 0 0 3
619 370
853 370
853 230
13 1 5 0 0 4224 0 10 7 0 0 3
619 379
929 379
929 258
14 1 6 0 0 8320 0 10 6 0 0 4
619 388
619 384
997 384
997 279
5 14 6 0 0 0 0 10 10 0 0 6
555 370
545 370
545 427
627 427
627 388
619 388
1 1 7 0 0 8320 0 1 10 0 0 4
403 236
478 236
478 316
555 316
1 4 2 0 0 8320 0 4 10 0 0 3
440 370
440 361
555 361
1 3 8 0 0 4224 0 2 10 0 0 4
422 309
504 309
504 343
555 343
1 0 9 0 0 4096 0 3 0 0 11 3
531 215
577 215
577 261
6 0 9 0 0 8320 0 10 0 0 11 4
549 388
535 388
535 306
549 306
7 2 9 0 0 0 0 10 10 0 0 6
619 316
623 316
623 261
549 261
549 334
555 334
10 1 2 0 0 0 0 10 5 0 0 5
619 343
680 343
680 283
694 283
694 291
9 1 2 0 0 0 0 10 5 0 0 5
619 334
680 334
680 283
694 283
694 291
8 1 2 0 0 0 0 10 5 0 0 5
619 325
680 325
680 283
694 283
694 291
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
263172 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.05 2
0
0 0 100 100 0 0
77 66 1487 276
0 0 0 0
1487 66
77 66
1487 66
1487 276
0 0
9.99575e-007 0 4.57143 4.14286 1e-006 1e-006
12409 0
0 3e-007 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
